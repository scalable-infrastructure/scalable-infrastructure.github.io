
<!DOCTYPE html>
<html lang="en">
  <head>
    <meta charset="utf-8">
    <title>Pages</title>
    
    <meta name="author" content="Andre Luckow">

    <!-- Le HTML5 shim, for IE6-8 support of HTML elements -->
    <!--[if lt IE 9]>
      <script src="http://html5shim.googlecode.com/svn/trunk/html5.js"></script>
    <![endif]-->

    <!-- Le styles -->
    <link href="/assets/themes/twitter/bootstrap/css/bootstrap.min.css" rel="stylesheet">
    <link href="/assets/themes/twitter/css/style.css?body=1" rel="stylesheet" type="text/css" media="all">

    <!-- Le fav and touch icons -->
  <!-- Update these with your own images
    <link rel="shortcut icon" href="images/favicon.ico">
    <link rel="apple-touch-icon" href="images/apple-touch-icon.png">
    <link rel="apple-touch-icon" sizes="72x72" href="images/apple-touch-icon-72x72.png">
    <link rel="apple-touch-icon" sizes="114x114" href="images/apple-touch-icon-114x114.png">
  -->
  </head>

  <body>

    <div class="navbar">
      <div class="navbar-inner">
        <div class="container">
          <a class="brand" href="/">Big Data und Large Scale Systems</a>
          <ul class="nav">
            
            
            


  
    
      
    
  
    
      
      	
      	<li><a href="/contact.html">Kontakt</a></li>
      	
      
    
  
    
      
    
  
    
      
      	
      	<li class="active"><a href="/pages.sv" class="active">Pages</a></li>
      	
      
    
  
    
      
    
  



          </ul>
        </div>
      </div>
    </div>

    <div class="container">

      <div class="content">
        
<div class="page-header">
  <!--h1>Pages </h1-->
  <h1>Pages </h1>
</div>

<div class="row">
  <div class="span12">
    

<h2>All Pages</h2>
<ul>




  
    
      
      	
      	<li><a href="/atom.xml">Atom Feed</a></li>
      	
      
    
  
    
      
      	
      	<li><a href="/contact.html">Kontakt</a></li>
      	
      
    
  
    
      
      	
      	<li><a href="/index.html">Überblick</a></li>
      	
      
    
  
    
      
      	
      	<li class="active"><a href="/pages.sv" class="active">Pages</a></li>
      	
      
    
  
    
      
      	
      	<li><a href="/sitemap.txt">Sitemap</a></li>
      	
      
    
  



</ul>

  </div>
</div>


      </div>

      <footer>
        <p>&copy; Andre Luckow 2012</p>
      </footer>

    </div> <!-- /container -->

    
  </body>
</html>

